module myfilter(
    input a,
    input b,
    input c,
    input d,
    output reg w,
    output reg x,
    output reg y,
    output reg z
);

// add your code here

endmodule
