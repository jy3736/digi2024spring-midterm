module shift_register(
    input wire clk,
    input wire rst,
    input wire L,        
    input wire r0,       
    input wire r1,       
    input wire r2,       
    output reg Q0,
    output reg Q1,
    output reg Q2
);

// add your code here

endmodule
