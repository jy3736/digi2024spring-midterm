module comb3i2o(
    input a,
    input b,
    input c,
    output reg x,
    output reg y
);

// add your code here

endmodule
